`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/12/2023 09:49:26 PM
// Design Name: 
// Module Name: tile_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tile_rom( 
        input [7:0]	  addr,
		output [7:0]  data );
		
		parameter ADDR_WIDTH = 8;
   parameter DATA_WIDTH =  8;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	// floor
	8'b10000011,
	8'b01100011,
	8'b01110000,
	8'b00010000,
	8'b00011000,
	8'b00001110,
	8'b00000010,
	8'b00000011,
	8'b10000011,
	8'b01100011,
	8'b01110000,
	8'b00010000,
	8'b00011000,
	8'b00001110,
	8'b00000010,
	8'b00000011,
	//wall
	8'b10000011,
	8'b01100011,
	8'b01110000,
	8'b00010000,
	8'b00011000,
	8'b00001110,
	8'b00000010,
	8'b00000011,
	8'b10000011,
	8'b01100011,
	8'b01110000,
	8'b00010000,
	8'b00011000,
	8'b00001110,
	8'b00000010,
	8'b00000011,
	//red door
	8'b11111111,
	8'b10100001,
	8'b10010001,
	8'b10100011,
	8'b11000101,
	8'b10001001,
	8'b10010001,
	8'b10001001,
	8'b11111111,
	8'b10100001,
	8'b10010001,
	8'b10100011,
	8'b11000101,
	8'b10001001,
	8'b10010001,
	8'b10001001,
	//blue door
	8'b11111111,
	8'b10100001,
	8'b10010001,
	8'b10100011,
	8'b11000101,
	8'b10001001,
	8'b10010001,
	8'b10001001,
	8'b11111111,
	8'b10100001,
	8'b10010001,
	8'b10100011,
	8'b11000101,
	8'b10001001,
	8'b10010001,
	8'b10001001,
	//lava
	8'b01000100,
	8'b00101000,
	8'b00010000,
	8'b00101000,
	8'b01000100,
	8'b10000010,
	8'b01000001,
	8'b00100010,
	8'b00010100,
	8'b00001000,
	8'b00001000,
	8'b00010100,
	8'b00100010,
	8'b01000001,
	8'b10000010,
	8'b01000100,
	//water
	8'b00000100,
	8'b00001010,
	8'b00000100,
	8'b00000000,
	8'b00100000,
	8'b01010000,
	8'b00100000,
	8'b00000000,
	8'b00000100,
	8'b00001010,
	8'b00000100,
	8'b00000000,
	8'b00100000,
	8'b01010000,
	8'b00100000,
	8'b00000000,
	//pressure plate
	8'b00000000,
	8'b00000000,
	8'b00011000,
	8'b00011000,
	8'b00011000,
	8'b00011000,
	8'b01111110,
	8'b01000010,
	8'b00100100,
	8'b00011000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b01111110,
	8'b10000001,
	8'b10000001,
	//puzzle door
	8'b11111111,
	8'b10000001,
	8'b10000001,
	8'b10000001,
	8'b10011001,
	8'b10100101,
	8'b10100101,
	8'b10011001,
	8'b10010001,
	8'b10011001,
	8'b10010001,
	8'b10011001,
	8'b10000001,
	8'b10000001,
	8'b10000001,
	8'b11111111,
	//level background
	8'b00010000,
	8'b00100000,
	8'b00010000,
	8'b00001000,
	8'b00010000,
	8'b00101000,
	8'b01000100,
	8'b00101000,
	8'b00010000,
	8'b00001000,
	8'b00000100,
	8'b00001000,
	8'b00010000,
	8'b00100000,
	8'b00010000,
	8'b00001000,
	//UNUSED
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	//UNUSED
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	//UNUSED
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	//UNUSED
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	//UNUSED
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	//UNUSED
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	//UNUSED
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000,
	8'b00000000
	};
		
	assign data = ROM[addr];	
	
endmodule

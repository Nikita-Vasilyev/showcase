`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/01/2023 08:36:39 PM
// Design Name: 
// Module Name: sprite_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sprite_rom(
        input [7:0]	  addr,
		output [63:0]  data );
		
    parameter ADDR_WIDTH = 8;
    parameter DATA_WIDTH =  64;
	logic [ADDR_WIDTH-1:0] addr_reg;
	
	// ROM definition, 2 bits color index for each pixel			
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	// fireboty stand
	// 0x0 = no color, 0x1 = black, 0x2 = light red, 0x3 = red, 0x4 = light yellow
	64'h0000000001000000,
    64'h0000100012101000,
    64'h0001210132212100,
    64'h0013231233232100,
    64'h0012323233332100,
    64'h0012323333333100,
    64'h0013333333333100,
    64'h0013313333133100,
    64'h0013141331413100,
    64'h0012313333133100,
    64'h0012333333332100,
    64'h0012333333332100,
    64'h0012313333332100,
    64'h0001331111321000,
    64'h0000133333310000,
    64'h0000011111100000,
    64'h0000001331000000,
    64'h0000013333100000,
    64'h0000133333310000,
    64'h0001333333331000,
    64'h0013333333333100,
    64'h0133113333113310,
    64'h0131013333101310,
    64'h0010013333100100,
    64'h0000013333100000,
    64'h0000013333100000,
    64'h0000133113310000,
    64'h0000131001310000,
    64'h0000131001310000,
    64'h0000131001310000,
    64'h0000131001310000,
    64'h0000111001110000,
    
    // fireboy right
    // 0x0 = no color, 0x1 = black, 0x2 = light red, 0x3 = red, 0x4 = light yellow
    64'h0001100000000000,
    64'h0013310000000000,
    64'h0112331000000000,
    64'h1231233100000000,
    64'h0123123310000000,
    64'h1313313311100000,
    64'h1231331333310000,
    64'h0123323333331000,
    64'h1312332331333100,
    64'h1231333314133100,
    64'h0133333331333100,
    64'h0123333333333100,
    64'h0012333133333100,
    64'h0001233311131000,
    64'h0000132223310000,
    64'h0000011111100000,
    64'h0000001331000000,
    64'h0000001331000000,
    64'h0000001331000000,
    64'h0000011331000000,
    64'h0000131333100000,
    64'h0001331333310000,
    64'h0013311331331000,
    64'h0013101331131000,
    64'h0001001331010000,
    64'h0000001331000000,
    64'h0000001331000000,
    64'h0000013331100000,
    64'h0000133313310000,
    64'h0001333101331000,
    64'h0001331000131000,
    64'h0000110000011000,
    
    // UNUSED (fireboy left)
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    
    // watergirl
    // 0x0 = no color, 0x1 = black, 0x2 = light blue, 0x3 = blue
    64'h0000001000000000,
    64'h0000013100000000,
    64'h0000132310000000,
    64'h0001113111110000,
    64'h0013321333321000,
    64'h0133231333233100,
    64'h1332331332333310,
    64'h1323313123333331,
    64'h0111133311111131,
    64'h0013313333133110,
    64'h0013121331213100,
    64'h0013333333333100,
    64'h0013333333133100,
    64'h0131331111231000,
    64'h0133133332210000,
    64'h1331011111100000,
    64'h1310001331000000,
    64'h0100013333100000,
    64'h0000133333310000,
    64'h0001333333331000,
    64'h0013333333333100,
    64'h0133113333113310,
    64'h0131013333101310,
    64'h0010013333100100,
    64'h0000013333100000,
    64'h0000013333100000,
    64'h0000133113310000,
    64'h0000131001310000,
    64'h0000131001310000,
    64'h0000131001310000,
    64'h0000131001310000,
    64'h0000111001110000,
    
    // watergirl right
    // 0x0 = no color, 0x1 = black, 0x2 = light blue, 0x3 = blue
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000011111010000,
    64'h0000133233131000,
    64'h0001332333133100,
    64'h0013323331333210,
    64'h0133233111332331,
    64'h1332311333123331,
    64'h1321133333311110,
    64'h1213333331333100,
    64'h1313323312133100,
    64'h1313232333333100,
    64'h1313323133333100,
    64'h1331333311131000,
    64'h1310133333310000,
    64'h0100011111100000,
    64'h0000001331000000,
    64'h0000001331000000,
    64'h0000001331000000,
    64'h0000011331000000,
    64'h0000131333100000,
    64'h0001331333310000,
    64'h0013311331331000,
    64'h0013101331131000,
    64'h0001001331010000,
    64'h0000001331000000,
    64'h0000001331000000,
    64'h0000013331100000,
    64'h0000133313310000,
    64'h0001333101331000,
    64'h0001331000131000,
    64'h0000110000011000,
    
    // UNUSED (watergirl left)
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    
    // UNUSED
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    
    // UNUSED
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000
    
	};
	
	assign data = ROM[addr];
    
endmodule
